module test

import math

const max_int = int(math.powi(2, 32))
