module html

pub type AttributeValue = string | bool
