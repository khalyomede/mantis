module css

type StyleBlock = Selector | Supports
