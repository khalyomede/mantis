module console

pub fn error(message string) {
    log(.error, message)
}
