module data

pub const internet_protocols = [
    "http"
    "https"
]
