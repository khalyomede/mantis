module console

pub struct Name {
    pub:
        name string
}
