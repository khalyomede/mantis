module cors

pub const default_headers = ["Content-Type", "Authorization", "Accept"]
