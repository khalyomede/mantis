module cors

pub const default_origins = ["*"]
