module console

pub struct Response {
    pub:
        output string
        code int
}
