module translation

pub enum Countable {
    zero
    one
    many
    any
}
