module console

pub fn info(message string) {
    log(.info, message)
}
