module data

pub const words = [
    "serendipity"
    "cascade"
    "luminous"
    "ephemeral"
    "mellifluous"
    "tranquil"
    "nebula"
    "pristine"
    "eloquent"
    "labyrinth"
    "whimsical"
    "ethereal"
]
