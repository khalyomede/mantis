module console

pub type ConsolePart = Program | Name | Argument | Flag | Opt
