module validation

pub type Value = string | int | u16 | u64 | i64
