module data

pub const person_last_names = [
    "Anderson"
    "Brown"
    "Smith"
]
