module data

pub const internet_top_level_domains = [
    "com"
    "io"
    "co.uk"
    "org"
]
