module data

pub const person_first_names = [
    "Adam"
    "John"
    "Mark"
];
