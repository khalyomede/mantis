module data

pub const company_names = [
    "Microsoft"
    "Apple"
    "Amazon"
    "Netflix"
    "Google"
    "Toyota"
    "Samsung"
    "Nike"
    "Coca-Cola"
    "Walmart"
    "Meta"
    "Sony"
    "Disney"
    "Nintendo"
    "Starbucks"
    "Adobe"
    "Intel"
    "Tesla"
    "BMW"
    "PayPal"
    "Spotify"
    "Twitter"
    "Airbnb"
    "Uber"
    "LinkedIn"
    "Nvidia"
    "Adidas"
    "Pepsi"
    "Honda"
    "FedEx"
    "Oracle"
    "Salesforce"
    "IBM"
    "Dell"
    "HP"
    "Cisco"
]
