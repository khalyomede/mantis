module css

pub type SelectorBlock = Rule | Selector
