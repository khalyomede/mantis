module translation

/**
 * @todo complete it
 */
pub enum Lang {
    en
    fr
    es
    cn
    ru
    ar
}
