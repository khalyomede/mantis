module cors

pub const default_max_age = 7200
