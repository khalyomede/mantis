module console

pub struct Program {
    pub:
        name string
}
