module generator

pub struct Country {
    pub:
        code CountryCode
}
