module http

pub enum SessionDriver {
    file
}
