module http

pub enum ServeMode {
    standalone
}
