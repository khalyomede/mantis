module database

pub enum DatabaseDriver {
    sqlite
}
