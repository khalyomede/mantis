module translation

pub enum Gender {
    feminine
    masculine
    neutral
}
