module console

pub fn debug(message string) {
    log(.debug, message)
}
