module console

type ConsolePart = Program | Name | Argument | Flag | Opt
