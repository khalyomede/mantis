module data

pub const internet_domains = [
  'gmail',
  'yahoo',
  'hotmail',
  'outlook',
  'proton',
  'example',
  'mail',
  'fastmail'
];
