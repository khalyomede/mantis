module data

pub const sentences = [
    "The meeting has been rescheduled."
    "Please review the attached document."
    "The project deadline is approaching."
    "We need to discuss the budget."
    "The client approved the proposal."
]
