module validation

pub type Value = string | int | u16
