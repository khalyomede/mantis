module console

type Part = Name | Argument | Flag | Opt
