module http

pub struct Middlewares {
    pub:
        before_route_match []Middleware
        after_route_match []Middleware
}
